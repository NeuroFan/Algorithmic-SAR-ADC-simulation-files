SRIVR10
*------------------ SRIVR-------------------           
*-------------------------------------------------

.subckt SRIVR10	SEL	D	CLK 	Pre	CLR	BI9	BI8	BI7	BI6	BI5	BI4	BI3	BI2	BI1	BI0	S9	S8	S7	S6	S5	S4	S3	S2	S1	S0

XMUX9	SEL	D	BI9	S9	Mux2-1 
XDFF9	S9	CLR	CLK	Pre	Q9	DFF

XMUX8	SEL	Q9	BI8	S8	Mux2-1 
XDFF8	S8	CLR	CLK	Pre	Q8	DFF

XMUX7	SEL	Q8	BI7	S7	Mux2-1 
XDFF7	S7	CLR	CLK	Pre	Q7	DFF

XMUX6	SEL	Q7	BI6	S6	Mux2-1 
XDFF6	S6	CLR	CLK	Pre	Q6	DFF

XMUX5	SEL	Q6	BI5	S5	Mux2-1 
XDFF5	S5	CLR	CLK	Pre	Q5	DFF

XMUX4	SEL	Q5	BI4	S4	Mux2-1 
XDFF4	S4	CLR	CLK	Pre	Q4	DFF

XMUX3	SEL	Q4	BI3	S3	Mux2-1 
XDFF3	S3	CLR	CLK	Pre	Q3	DFF

XMUX2	SEL	Q3	BI2	S2	Mux2-1 
XDFF2	S2	CLR	CLK	Pre	Q2	DFF

XMUX1	SEL	Q2	BI1	S1	Mux2-1 
XDFF1	S1	CLR	CLK	Pre	Q1	DFF

XMUX0	SEL	Q1	BI0	S0	Mux2-1 
XDFF0	S0	CLR	CLK	Pre	Q0	DFF

.ends  SRIVR10 


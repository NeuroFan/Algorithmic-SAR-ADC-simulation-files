*-------------------------------------------------
*------------------ NOR8-------------------           
*-------------------------------------------------

.subckt NOR8	I1	I2	I3	I4	I5	I6	I7	I8	Out 

XR4-1	I1	I2	I3	I4	X1	OR4 
XR4-2	I5	I6	I7	I8	X2	OR4 

XNOR	X1	X2	Out	NOR2 


.ends  NOR8 

*-------------------------------------------------
*----------------------NOT------------------------           
*-------------------------------------------------

.subckt NOT  iin   oin
Mni1	oin      iin      ss	ss	N_10_SP	W=125n	L=0.09u	M=2    
Mpi1	oin      iin      ddd	ddd	P_10_SP	W=250n	L=0.09u	M=2   
.ends  NOT 
*-------------------------------------------------
*----------------------NOTD------------------------           
*-------------------------------------------------

.subckt NOTD  In   Out
Mni1	Out      In      ss	ss	N_10_SP	W=500n	L=0.09u	M=2    
Mpi1	Out      In      dd	dd	P_10_SP	W=1u	L=0.09u	M=2   
.ends  NOTD 
*-------------------------------------------------
*------------------ AND4-------------------           
*-------------------------------------------------

.subckt AND4	I1	I2	I3	I4	Out 

XAND1	I1	I2	X1	AND2 
XAND2	I3	I4	X2	AND2 

XAND	X1	X2	Out	AND2 


.ends  AND4 

*-------------------------------------------------
*------------------ ADSBN-------------------           
*-------------------------------------------------

.subckt ADSBN	B0	BD0	B1	BD1	B2	BD2	B3	BD3	B4	BD4
+B5	BD5	B6	BD6	B7	BD7	SB0	SB1	SB2	SB3	SB4
+SB5	SB6	SB7	SB8	SB9


XXOR0	B9	BD9	SB9	XOR_4ND

XXOR1	B8	BD8	X9	XOR_4ND
XNOT0	SB9	SBN9	NOT
XAND0	X9	SBN9	SB8	AND2

XXOR2	B7	BD7	X8	XOR_4ND
XOR1	SB9	SB8	O9	OR2
XNOT1	O9	OB9	NOT
XAND1	OB9	X8	SB7	AND2

XXOR3	B6	BD6	X7	XOR_4ND
XOR2	O9	SB7	O8	OR2
XNOT2	O8	OB8	NOT
XAND2	OB8	X7	SB6	AND2

XXOR4	B5	BD5	X6	XOR_4ND
XOR3	O8	SB6	O7	OR2
XNOT3	O7	OB7	NOT
XAND3	OB7	X6	SB5	AND2

XXOR5	B4	BD4	X5	XOR_4ND
XOR4	O7	SB5	O6	OR2
XNOT4	O6	OB6	NOT
XAND4	OB6	X5	SB4	AND2

XXOR6	B3	BD3	X4	XOR_4ND
XOR5	O6	SB4	O5	OR2
XNOT5	O5	OB5	NOT
XAND5	OB5	X4	SB3	AND2

XXOR7	B2	BD2	X3	XOR_4ND
XOR6	O5	SB3	O4	OR2
XNOT6	O4	OB4	NOT
XAND6	OB4	X3	SB2	AND2

XOR7	O4	SB2	O3	OR2
XNOT7	O3	OB3	NOT
XAND7	OB3	DD	SB1	AND2


XOR8	O3	SB1	O2	OR2
XNOT8	O2	OB2	NOT
XAND8	OB2	DD	SB0	AND2


.ends  ADSBN 

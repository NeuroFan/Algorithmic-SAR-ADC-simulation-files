*-------------------------------------------------
*------------------ ADSB-------------------           
*-------------------------------------------------

.subckt ADSB	B0	BD0	B1	BD1	B2	BD2	B3	BD3	B4	BD4
+B5	BD5	B6	BD6	B7	BD7	SB0	SB1	SB2	SB3	SB4
+SB5	SB6	SB7	SB8	SB9


XXOR0	B0	BD0	SB0	XOR_4ND

XXOR1	B1	BD1	X1	XOR_4ND
XNOT0	SB0	SBN0	NOT
XAND0	X1	SBN0	SB1	AND2

XXOR2	B2	BD2	X2	XOR_4ND
XOR1	SB0	SB1	O0	OR2
XNOT1	O0	OB0	NOT
XAND1	OB0	X2	SB2	AND2

XXOR3	B3	BD3	X3	XOR_4ND
XOR2	O0	SB2	O1	OR2
XNOT2	O1	OB1	NOT
XAND2	OB1	X3	SB3	AND2

XXOR4	B4	BD4	X4	XOR_4ND
XOR3	O1	SB3	O2	OR2
XNOT3	O2	OB2	NOT
XAND3	OB2	X4	SB4	AND2

XXOR5	B5	BD5	X5	XOR_4ND
XOR4	O2	SB4	O3	OR2
XNOT4	O3	OB3	NOT
XAND4	OB3	X5	SB5	AND2

XXOR6	B6	BD6	X6	XOR_4ND
XOR5	O3	SB5	O4	OR2
XNOT5	O4	OB4	NOT
XAND5	OB4	X6	SB6	AND2

XXOR7	B7	BD7	X7	XOR_4ND
XOR6	O4	SB6	O5	OR2
XNOT6	O5	OB5	NOT
XAND6	OB5	X7	SB7	AND2

XOR7	O5	SB7	O6	OR2
XNOT7	O6	OB6	NOT
XAND7	OB6	DD	SB8	AND2


XOR8	O6	SB8	O7	OR2
XNOT8	O7	OB7	NOT
XAND8	OB7	DD	SB9	AND2


.ends  ADSB 
